module LAC(c, gout, pout, Cin, g, p);
      output[1:0] c;
      output gout, pout;
      input Cin;
      input[1:0] g, p;

      assign c[0] = Cin;
      assign c[1] = g[0] | (p[0] & Cin);
      assign gout = g[1] | (p[1] & g[0]);
      assign pout = p[1] & p[0];
endmodule
